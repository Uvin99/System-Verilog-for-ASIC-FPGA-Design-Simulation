module n_adder #(
    parameter N=4
)(
    inpiut logic signed
);









endmodule